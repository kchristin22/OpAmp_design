** Profile: "SCHEMATIC1-ACsweep"  [ C:\Users\chris\Documents\spice\miller_op_amp_9994-PSpiceFiles\SCHEMATIC1\ACsweep.sim ] 

** Creating circuit file "ACsweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../miller_op_amp_9994-pspicefiles/miller_op_amp_9994.lib" 
* From [PSPICE NETLIST] section of C:\SPB_DATA\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 40 1 1e+10
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
