** Profile: "SCHEMATIC1-R_sweep"  [ c:\users\chris\documents\spice\miller_op_amp_9994-PSpiceFiles\SCHEMATIC1\R_sweep.sim ] 

** Creating circuit file "R_sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../miller_op_amp_9994-pspicefiles/miller_op_amp_9994.lib" 
* From [PSPICE NETLIST] section of C:\SPB_DATA\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.STEP LIN PARAM RVAL 100 110 2 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
